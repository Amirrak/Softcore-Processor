library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity registre is
    port (
        dataIn          : in std_logic_vector(7 downto 0);  -- entree donnee sur 8 bits
        cs, rst, clk    : in std_logic;                     -- chip select, reset, et clock
        q               : out std_logic_vector(7 downto 0)  -- sortie du registre sur 8 bits
    );
end registre;

architecture Behavioral of registre is

begin
    
    process(clk)
    begin
    
        if (clk'event and clk='1') then
            if rst = '1' then
                q <= (others => '0');
            else
                if cs = '1' then
                    q <= dataIn;
                end if;
            end if;
        end if;
        
    end process;

end Behavioral;
